// Copyright 2017 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the “License”); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

module boot_code_latch
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:838] [31:0] mem = {
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h00000013,
32'h0100006f,
32'h0100006f,
32'h0080006f,
32'h0040006f,
32'h0000006f,
32'h00000093,
32'h81868106,
32'h82868206,
32'h83868306,
32'h84868406,
32'h85868506,
32'h86868606,
32'h87868706,
32'h88868806,
32'h89868906,
32'h8a868a06,
32'h8b868b06,
32'h8c868c06,
32'h8d868d06,
32'h8e868e06,
32'h8f868f06,
32'h00100117,
32'hf3010113,
32'h00001d17,
32'hc48d0d13,
32'h00001d97,
32'hc40d8d93,
32'h01bd5763,
32'h000d2023,
32'hdde30d11,
32'h0513ffad,
32'h05930000,
32'h00ef0000,
32'h11012180,
32'h1000ce22,
32'h07a387aa,
32'h4783fef4,
32'h0733fef4,
32'h07b700f0,
32'h07d11a10,
32'hf793439c,
32'hdbf50207,
32'h1a1007b7,
32'h07d1c398,
32'h77134398,
32'hdf6d0407,
32'h44720001,
32'h80826105,
32'hce061101,
32'h1000cc22,
32'h242387aa,
32'h8736feb4,
32'hfef407a3,
32'h072387b2,
32'h87bafef4,
32'hfef406a3,
32'hfef44783,
32'hfe842703,
32'hfee44683,
32'h45a1863a,
32'h00ef853e,
32'h47830c90,
32'h4581fed4,
32'h00ef853e,
32'h2a951bd0,
32'h40f20001,
32'h61054462,
32'h71798082,
32'hd422d606,
32'h87aa1800,
32'hfcf40fa3,
32'h46014681,
32'h451545a1,
32'h097000ef,
32'h00ef4521,
32'h458114d0,
32'h00ef4501,
32'h47831110,
32'h4581fdf4,
32'h00ef853e,
32'h2a1517d0,
32'hfef40793,
32'h853e45a1,
32'h249000ef,
32'hfef44783,
32'hf3f98b85,
32'h50b20001,
32'h61455422,
32'h11018082,
32'hcc22ce06,
32'h26231000,
32'h2423fea4,
32'h2223feb4,
32'h2783fec4,
32'h07a2fec4,
32'h02000693,
32'h45a1863e,
32'h0eb00513,
32'h033000ef,
32'hfe842503,
32'h0e7000ef,
32'h45114581,
32'h0ab000ef,
32'h45094581,
32'h11b000ef,
32'hfe842583,
32'hfe442503,
32'h1e9000ef,
32'h40f20001,
32'h61054462,
32'h11018082,
32'hcc22ce06,
32'h26231000,
32'h2423fea4,
32'h2223feb4,
32'h468dfec4,
32'h45814601,
32'h35ed4519,
32'hfec42783,
32'h863e46e1,
32'h450945a1,
32'h7d6000ef,
32'hfe842783,
32'h00ef853e,
32'h45810890,
32'h00ef450d,
32'h27830c50,
32'h85befe84,
32'hfe442503,
32'h115000ef,
32'h450920bd,
32'h00013709,
32'h446240f2,
32'h80826105,
32'hd6067179,
32'h1800d422,
32'hfca42e23,
32'hfcb42c23,
32'hfe042623,
32'h468da815,
32'h45814601,
32'h35694519,
32'h4661468d,
32'hfdc42583,
32'h0d700513,
32'h45093db5,
32'h270335d9,
32'h6785fdc4,
32'h2e2397ba,
32'h2783fcf4,
32'h0785fec4,
32'hfef42623,
32'hfec42703,
32'hfd842783,
32'hfcf763e3,
32'h50b20001,
32'h61455422,
32'h11418082,
32'hc422c606,
32'h00010800,
32'h07d000ef,
32'hf71387aa,
32'h478503f7,
32'hfef71ae3,
32'h40b20001,
32'h01414422,
32'h11018082,
32'hcc22ce06,
32'ha7b71000,
32'h07911a10,
32'ha7b74398,
32'h07911a10,
32'h00876713,
32'ha7b7c398,
32'h07911a10,
32'ha7b74398,
32'h07911a10,
32'h00276713,
32'ha7b7c398,
32'h07911a10,
32'ha7b74398,
32'h07911a10,
32'h01076713,
32'h2623c398,
32'ha039fe04,
32'h27830001,
32'h0785fec4,
32'hfef42623,
32'hfec42703,
32'h87936785,
32'hd5e395f7,
32'h47fdfee7,
32'ha7b7873e,
32'h07911a10,
32'h0007a283,
32'h0022e293,
32'h0057a023,
32'h1a1007b7,
32'ha28307b1,
32'hf2930007,
32'he2b30c02,
32'ha02300e2,
32'h478d0057,
32'h07b7873e,
32'h07b11a10,
32'h0007a283,
32'h0802e293,
32'h0057a023,
32'h1a100837,
32'h00e82023,
32'h08118321,
32'h00e82023,
32'h07f2f293,
32'h0057a023,
32'h0a700793,
32'h07b7873e,
32'h07b11a10,
32'h0007a283,
32'h0802e293,
32'h0057a023,
32'h1a100837,
32'h23030821,
32'h73130008,
32'h63330183,
32'h202300e3,
32'hf2930068,
32'ha02307f2,
32'h479d0057,
32'h0ff7f713,
32'h1a1037b7,
32'hc3980791,
32'h45054585,
32'h06f000ef,
32'h82be4785,
32'h27b74305,
32'ha3831a10,
32'h13330007,
32'h43130053,
32'hf3b3fff3,
32'ha0230063,
32'h46850077,
32'h45814601,
32'h39dd4519,
32'h46214685,
32'h04200593,
32'h31ed4505,
32'h3b154501,
32'h46014685,
32'h05134581,
32'h39e90350,
32'h873e4785,
32'h1a1027b7,
32'ha2830791,
32'hd2b30007,
32'hf29300e2,
32'h87960012,
32'hfef405a3,
32'hfeb44783,
32'h4705c789,
32'h00e78563,
32'h2295a029,
32'h2cc1a019,
32'ha0010001,
32'h2e237129,
32'h2c231211,
32'h02801281,
32'heca42623,
32'hecb42423,
32'hecc42223,
32'h10000793,
32'hfef42623,
32'hed840793,
32'hfcf42c23,
32'hfe0405a3,
32'hec442703,
32'h0ff00793,
32'h00e7e663,
32'hec442783,
32'hfef42623,
32'hfe042223,
32'h0001a8e5,
32'h003000ef,
32'h873e87aa,
32'h05300793,
32'hfef71ae3,
32'hfe042023,
32'h00efa00d,
32'h87aa7ec0,
32'h2783873e,
32'h0693fe04,
32'h97b6ff04,
32'heee78423,
32'hfe042783,
32'h20230785,
32'h2783fef4,
32'h2703fe04,
32'hece3fec4,
32'h2703fce7,
32'h0793fec4,
32'h0e631000,
32'h278300f7,
32'hf793fec4,
32'h8b8d0ff7,
32'h0ff7f793,
32'h07b34711,
32'h05a340f7,
32'h2e23fef4,
32'ha005fc04,
32'hfdc42703,
32'hfec42783,
32'h071397ba,
32'h97baff04,
32'hee078423,
32'hfdc42783,
32'h2e230785,
32'h4783fcf4,
32'h2703feb4,
32'h4de3fdc4,
32'h4783fcf7,
32'h2703feb4,
32'h97bafec4,
32'hfef42623,
32'h02000513,
32'h27833ead,
32'h9713fe44,
32'h27830087,
32'h973eec84,
32'hfec42783,
32'h0693078e,
32'h8636ed84,
32'h853a85be,
32'h27833179,
32'h0785fe44,
32'h270307a2,
32'h07b3ec44,
32'h071340f7,
32'h74631000,
32'h079300f7,
32'h26231000,
32'h2783fef4,
32'h0785fe44,
32'hfef42223,
32'hfe442703,
32'hecc42783,
32'hf0f761e3,
32'hfd842783,
32'h2083853e,
32'h240313c1,
32'h61311381,
32'h71398082,
32'hdc22de06,
32'h45410080,
32'h00013619,
32'h6e2000ef,
32'hffed87aa,
32'hfd040793,
32'h0593863e,
32'h45110200,
32'h079336e9,
32'h863efc84,
32'h02000593,
32'h3e754561,
32'hfcc40793,
32'h0593863e,
32'h45410200,
32'h2703367d,
32'h57fdfc84,
32'h00f70763,
32'hfd042703,
32'h106357fd,
32'h468d02f7,
32'h45814601,
32'h34fd4519,
32'h4601468d,
32'h05134581,
32'h34cd0600,
32'h36354509,
32'h2783a091,
32'h8793fd04,
32'h28231007,
32'h2703fcf4,
32'h6785fd04,
32'h8ff917fd,
32'h2783c791,
32'h83b1fd04,
32'ha0210785,
32'hfd042783,
32'h262383b1,
32'h2783fef4,
32'h2703fcc4,
32'h85bafc84,
32'h3eed853e,
32'hfec42583,
32'h3ecd4501,
32'h3cb14545,
32'h02800613,
32'h45054581,
32'h242333e5,
32'h454dfea4,
32'h278334a9,
32'h439cfe84,
32'hfef42223,
32'hfe842783,
32'h282343dc,
32'h2783fcf4,
32'h539cfe84,
32'hfef42023,
32'hfe842783,
32'h26234b9c,
32'h2783fcf4,
32'h4bdcfe84,
32'hfcf42e23,
32'hfe842783,
32'h2c2353dc,
32'h2783fcf4,
32'h863efd04,
32'hfe442583,
32'hfe042503,
32'h45513b51,
32'h27833aed,
32'h2603fcc4,
32'h85befdc4,
32'hfd842503,
32'h45553341,
32'h23d132dd,
32'h0ba387aa,
32'h4703fcf4,
32'h47d9fd74,
32'h02f71063,
32'hfd042783,
32'h250385be,
32'h2af5fe44,
32'hfcc42783,
32'hfdc42583,
32'h2ac5853e,
32'ha0392829,
32'hfd744703,
32'h136347dd,
32'h203100f7,
32'h50f20001,
32'h61215462,
32'h71398082,
32'hdc22de06,
32'h07930080,
32'h863efc84,
32'h10000593,
32'h34a54501,
32'hfd442783,
32'hfef42623,
32'hfe442783,
32'hfef42423,
32'hfc842783,
32'h2783873e,
32'h85befd04,
32'hfcc42783,
32'hfec42683,
32'h853a863e,
32'h2783280d,
32'h873efd84,
32'hfe042783,
32'h278385be,
32'h2683fdc4,
32'h863efe84,
32'h2821853a,
32'hfd442783,
32'h08078793,
32'h00078067,
32'h50f20001,
32'h61215462,
32'h71798082,
32'hd422d606,
32'h2e231800,
32'h2c23fca4,
32'h2a23fcb4,
32'h2823fcc4,
32'h6785fcd4,
32'hfef42623,
32'hfd442783,
32'h00478693,
32'hfd442703,
32'h41f75793,
32'h973e83f9,
32'h07b38b0d,
32'h87b340f7,
32'h2a2340f6,
32'h2703fcf4,
32'h6785fd44,
32'h00f75663,
32'hfd442783,
32'hfef42623,
32'hfe042423,
32'h2783a889,
32'h078efec4,
32'hfd042603,
32'h250385be,
32'h3255fdc4,
32'hfe842783,
32'h07b20785,
32'hfd442703,
32'h40f707b3,
32'h53636705,
32'h678500f7,
32'hfef42623,
32'hfd042703,
32'h97ba6785,
32'hfcf42823,
32'hfdc42703,
32'h97ba6785,
32'hfcf42e23,
32'hfe842783,
32'h24230785,
32'h2703fef4,
32'h2783fe84,
32'h44e3fd84,
32'h34b5faf7,
32'h50b20001,
32'h61455422,
32'h71798082,
32'h1800d622,
32'hfca42e23,
32'h873287ae,
32'hfcf40da3,
32'h0d2387ba,
32'h2623fcf4,
32'ha885fe04,
32'hfec42783,
32'hfdc42703,
32'hc78397ba,
32'h05a30007,
32'h2223fef4,
32'ha091fe04,
32'hfda44783,
32'h01a38b85,
32'h4783fef4,
32'h8385fda4,
32'hfcf40d23,
32'hfe344703,
32'hfeb44783,
32'h08638b85,
32'h478300f7,
32'hc793fda4,
32'h0d23f8c7,
32'h4783fcf4,
32'h8385feb4,
32'hfef405a3,
32'hfe442783,
32'h22230785,
32'h2703fef4,
32'h479dfe44,
32'hfae7dce3,
32'hfec42783,
32'h26230785,
32'h4783fef4,
32'h2703fdb4,
32'h45e3fec4,
32'h4783f8f7,
32'h853efda4,
32'h61455432,
32'h71398082,
32'hdc22de06,
32'h26230080,
32'h2423fca4,
32'h07a3fcb4,
32'h2783fe04,
32'h8389fc84,
32'hfef42023,
32'hfe042423,
32'h2783a0a1,
32'h0713fcc4,
32'h863afdc4,
32'h02000593,
32'h3895853e,
32'hfcc42783,
32'h26230791,
32'h2783fcf4,
32'h17f1fc84,
32'hfcf42423,
32'hfef44703,
32'hfdc40793,
32'h4591863a,
32'h3711853e,
32'h07a387aa,
32'h2783fef4,
32'h0785fe84,
32'hfef42423,
32'hfe842783,
32'hfe042703,
32'hfae7e9e3,
32'hfc042c23,
32'hfc842783,
32'h2783c7bd,
32'h0713fcc4,
32'h863afdc4,
32'h02000593,
32'h3821853e,
32'hfe042223,
32'h2783a035,
32'h078efe44,
32'h0ff00713,
32'h00f717b3,
32'h2783873e,
32'h8f7dfdc4,
32'hfd842783,
32'h2c2397ba,
32'h2783fcf4,
32'h0785fe44,
32'hfef42223,
32'hfe442783,
32'hfc842703,
32'hfce7e7e3,
32'hfc842783,
32'h0ff7f713,
32'hfef44683,
32'hfd840793,
32'h85ba8636,
32'h3da5853e,
32'h07a387aa,
32'h4783fef4,
32'h853efef4,
32'hedaff0ef,
32'h50f20001,
32'h61215462,
32'h71798082,
32'h1800d622,
32'hfca42e23,
32'hfcb42c23,
32'hfcc42a23,
32'hfcd42823,
32'h02000713,
32'hfd842783,
32'h40f707b3,
32'hfdc42703,
32'h00f717b3,
32'hfef42623,
32'h02000713,
32'hfd042783,
32'h40f707b3,
32'hfd442703,
32'h00f717b3,
32'hfef42423,
32'h1a1037b7,
32'h270307a1,
32'hc398fec4,
32'h1a1037b7,
32'h270307b1,
32'hc398fe84,
32'hfd842783,
32'h03f7f693,
32'hfd042783,
32'h00879713,
32'h87936791,
32'h8f7df007,
32'h1a1037b7,
32'h8f5507c1,
32'h0001c398,
32'h61455432,
32'h11018082,
32'h1000ce22,
32'hfea42623,
32'hfeb42423,
32'hfe842783,
32'h86be07c2,
32'hfec42703,
32'h17fd67c1,
32'he7338ff9,
32'h37b700f6,
32'h07d11a10,
32'h0001c398,
32'h61054472,
32'h71798082,
32'h1800d622,
32'hfca42e23,
32'h1a1037b7,
32'h439c07c1,
32'hfef42623,
32'hfdc42783,
32'h873e07c2,
32'hfec42783,
32'h67c186be,
32'h8ff517fd,
32'h26238fd9,
32'h37b7fef4,
32'h07c11a10,
32'hfec42703,
32'h0001c398,
32'h61455432,
32'h11018082,
32'h1000ce22,
32'hfea42623,
32'hfeb42423,
32'hfe842783,
32'h470507a1,
32'h00f71733,
32'h87936785,
32'h76b3f007,
32'h470500f7,
32'hfec42783,
32'h00f717b3,
32'h0ff7f713,
32'h1a1037b7,
32'hc3988f55,
32'h44720001,
32'h80826105,
32'hce221101,
32'h37b71000,
32'h439c1a10,
32'hfef42623,
32'hfec42783,
32'h4472853e,
32'h80826105,
32'hd6227179,
32'h2e231800,
32'h2c23fca4,
32'h2783fcb4,
32'h8795fd84,
32'h7ff7f793,
32'hfef42623,
32'hfd842783,
32'hc7918bfd,
32'hfec42783,
32'h26230785,
32'h2423fef4,
32'ha81dfe04,
32'h37b70001,
32'h439c1a10,
32'hf71387e1,
32'h479d0ff7,
32'hfee7c9e3,
32'hfe842783,
32'h2703078a,
32'h973efdc4,
32'h1a1037b7,
32'h431807e1,
32'h2783c398,
32'h0785fe84,
32'hfef42423,
32'hfe842703,
32'hfec42783,
32'hfcf742e3,
32'h54320001,
32'h80826145,
32'hd6227179,
32'h2e231800,
32'h2c23fca4,
32'h2783fcb4,
32'h8795fd84,
32'h7ff7f793,
32'hfef42623,
32'hfd842783,
32'hc7918bfd,
32'hfec42783,
32'h26230785,
32'h2423fef4,
32'ha815fe04,
32'h37b70001,
32'h439c1a10,
32'hf79387c1,
32'hdbf50ff7,
32'h1a1037b7,
32'h02078713,
32'hfe842783,
32'h2683078a,
32'h97b6fdc4,
32'hc3984318,
32'hfe842783,
32'h24230785,
32'h2703fef4,
32'h2783fe84,
32'h43e3fec4,
32'h0001fcf7,
32'h61455432,
32'h71798082,
32'h1800d622,
32'hfca42e23,
32'hfcb42c23,
32'h1a10a7b7,
32'h2623439c,
32'h4705fef4,
32'hfdc42783,
32'h00f717b3,
32'hfff7c713,
32'hfec42783,
32'h26238ff9,
32'h2703fef4,
32'h2783fd84,
32'h1733fdc4,
32'h278300f7,
32'h8fd9fec4,
32'hfef42623,
32'h1a10a7b7,
32'hfec42703,
32'h0001c398,
32'h61455432,
32'h11418082,
32'h0800c622,
32'h07b70001,
32'h07d11a10,
32'hf713439c,
32'h47850017,
32'hfef719e3,
32'h1a1007b7,
32'hf793439c,
32'h853e0ff7,
32'h01414432,
32'h00008082,
32'h00000000,
32'h00000000,
32'h00000000};

  logic [9:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule